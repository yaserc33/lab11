class c_145_4;
    int j = 4;
    rand bit[1:0] addr; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (yapp_tx_seqs.sv:126)
    {
       (addr == j);
    }
endclass

program p_145_4;
    c_145_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxxz0101zxz1x1xz10001010z0xx00zzxzxzzxzxzxzzzxxzzzxxzxzzzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
