class c_66_4;
    int j = 4;
    rand bit[1:0] addr; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (yapp_tx_seqs.sv:126)
    {
       (addr == j);
    }
endclass

program p_66_4;
    c_66_4 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zzz0zzz1100zxx1x0z1zx1zz11101xzzzxzxxxxxxxzzzxxxxxxzzxxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
