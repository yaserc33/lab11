class c_165_1;
    int i = 21;
    rand bit[5:0] length; // rand_mode = ON 

    constraint length2_this    // (constraint_mode = ON) (../sv/yapp_packet.sv:78)
    {
       (length < 6'hf);
    }
    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (yapp_tx_seqs.sv:126)
    {
       (length == i);
    }
endclass

program p_165_1;
    c_165_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx0xx1z0z0z01zxzx0101z0z0z0zz10xzzzxzzxxzxxzzzxzzxxzxxzxzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
